module TB_HitMissLogic();
logic [35:0] tagAddress,tagBloque1,tagBloque2,tagBloque3,tagBloque4;
logic vBit1,vBit2,vBit3,vBit4;
logic hit;

HitMissLogic dut(tagAddress,tagBloque1,tagBloque2,tagBloque3,tagBloque4,vBit1,vBit2,vBit3,vBit4,hit);

initial begin
tagAddress=36'b000000000000000000000000010000000000;
tagBloque1=36'b000000000000000000000000000000000000;
tagBloque2=36'b110000000000000000000000000000000000;
tagBloque3=36'b000000000000000000000000010000000000;
tagBloque4=36'b000000000100000000100000000000000000;
vBit1=1;vBit2=1;vBit3=1;vBit4=1; #10;
tagAddress=36'b000000000000000000000000010000000000;
tagBloque1=36'b000000000000000000000000000000000000;
tagBloque2=36'b110000000000000000000000000000000000;
tagBloque3=36'b000000000000000000000000000000000100;
tagBloque4=36'b000000000100000000100000000000000000;
vBit1=1;vBit2=1;vBit3=1;vBit4=1; #10;
tagAddress=36'b000000000000000000000000000000000001;
tagBloque1=36'b000000000000000000000000000000000000;
tagBloque2=36'b110000000000000000000000000000000000;
tagBloque3=36'b000000000000000000000000000000000100;
tagBloque4=36'b000000000000000000000000000000000000;
vBit1=1;vBit2=1;vBit3=1;vBit4=1; #10;
tagAddress=36'b000000000000000000000000000000000001;
tagBloque1=36'b000000000000000000000000000000000000;
tagBloque2=36'b110000000000000000000000000000000000;
tagBloque3=36'b000000000000000000000000000000000100;
tagBloque4=36'b000000000000000000000000000000000001;
vBit1=1;vBit2=1;vBit3=1;vBit4=1; #10;

end

endmodule